simple_circuit1
R1 n1 n2 1
R2 n2 n3 1
R3 n3 n4 1
V1 n1 0 4
I1 n4 0 1
.print dc v(*)
.op
.end